grammar custom:host:abstractsyntax;


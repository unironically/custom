grammar custom:host:typing;

imports custom:host:abstractsyntax;

aspect production file
top::File ::= ds::TopDecls
{
}
grammar custom:host:abstractsyntax;

nonterminal File with location;

abstract production file
top::File ::= ds::TopDecls
{}